Library ieee;
use ieee.std_logic_1164.all;
LIBRARY altera_mf;
USE lpm.lpm_components.all;